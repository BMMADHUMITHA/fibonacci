`include "design.v"
`include "fib_trans.sv"
`include "fib_gen.sv"
`include "fib_intf.sv"
`include "fib_bfm.sv"
`include "fib_env.sv"
`include "fib_test.sv"
`include "tb_fib_top.sv"





